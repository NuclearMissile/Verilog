`timescale 1ns / 1ps

module RSA(
    
);

endmodule // RSA